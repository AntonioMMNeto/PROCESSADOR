module UControle(IP_endereco,RET_endereco,IR_opcode,MAR_saida,TOS_saida,Dados);
