`timescale 10ns/1ns
module tb_Barramento;


parameter Largura_barramento=16;

reg [Largura_barramento-1:0]io_tb[3:0];
wire [Largura_barramento-1:0]io_out_tb[5:4];
reg [1:0] ctrl_tb[5:0]; //bit 0 ler; bit 1 escrever
reg clk_tb;
reg [Largura_barramento-1:0] io_in_tb;




Barramento barramento_tb (.io_0(io_tb[0]),.io_1(io_tb[1]),.io_2(io_tb[2]),.io_3(io_tb[3]),.io_4(io_out_tb[4]),.io_5(io_out_tb[5]),.ctrl_0(ctrl_tb[0]),.ctrl_1(ctrl_tb[1]),.ctrl_2(ctrl_tb[2]),.ctrl_3(ctrl_tb[3]),.ctrl_4(ctrl_tb[4]),.ctrl_5(ctrl_tb[5]),.clk(clk_tb));

/*assign io_tb[0]=io_in_tb[0];
assign io_tb[1]=io_in_tb[1];
assign io_tb[2]=io_in_tb[2];
assign io_tb[3]=io_in_tb[3];
assign io_tb[4]=io_in_tb[4];
assign io_tb[5]=io_in_tb[5];*/

integer x,y;
always
begin
	for(x=0;x<4;x=x+1)
	begin
		for(y=4;y<5;y=y+1)
			begin
					ctrl_tb[x]=2'b10;
					ctrl_tb[y]=2'b01;
					#10 clk_tb=1;
					#10 io_tb[x]=2;
					$monitor("Valor de sa�da na Porta %d :%d",y,io_out_tb[y]);
					#10 clk_tb=0;
			end
	end
end
endmodule
